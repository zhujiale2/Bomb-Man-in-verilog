`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:33:41 01/06/2014 
// Design Name: 
// Module Name:    winmap 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module winmap(	
	input wire clk,
	input wire [9:0] px, py,
	output wire end_on
);
	reg out;
	reg [1:160] map [1:120];
	initial begin
      map[120] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[119] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[118] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[117] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[116] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[115] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[114] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[113] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[112] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[111] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[110] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[109] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[108] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[107] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[106] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[105] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[104] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[103] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[102] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[101] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[100] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[99] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[98] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[97] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[96] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[95] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[94] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[93] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[92] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[91] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[90] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[89] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[88] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[87] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[86] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[85] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[84] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[83] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[82] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[81] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[80] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[79] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[78] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[77] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[76] = 160'b00000000000001111111100000000000000111111110000000000000000000000000001111111111111000000000000000000011111110000000000000000111111110000000;
      map[75] = 160'b00000000000001111111110000000000000111111111000000000000000000000000001111111111111000000000000000000011111110000000000000001111111110000000;
      map[74] = 160'b00000000000001111111110000000000000111111111000000000000000000000000001111111111111000000000000000000011111110000000000000001111111110000000;
      map[73] = 160'b00000000000001111111110000000000000111111111000000000000000000000000001111111111111000000000000000000011111110000000000000011111111110000000;
      map[72] = 160'b00000000000011111111110000000000001111111111100000000000000000000000001111111111111000000000000000000011111110000000000000011111111110000000;
      map[71] = 160'b00000000000011111111111000000000001111111111100000000000000000000000001111111111111000000000000000000011111110000000000000111111111110000000;
      map[70] = 160'b00000000000011111111111000000000001111111111100000000000000000000000001111111111111000000000000000000011111110000000000001111111111110000000;
      map[69] = 160'b00000000000011111111111000000000001111111111100000000000000000000000000011111111000000000000000000000011111110000000000001111111111110000000;
      map[68] = 160'b00000000000111111111111100000000011111111111110000000000000000000000000011111111000000000000000000000011111110000000000011111111111110000000;
      map[67] = 160'b00000000000111111111111100000000011111111111110000000000000000000000000011111111000000000000000000000011111110000000000111111111111110000000;
      map[66] = 160'b00000000000111111111111100000000011111111111110000000000000000000000000011111111000000000000000000000011111110000000000111111111111110000000;
      map[65] = 160'b00000000000111111111111100000000011111101111110000000000000000000000000011111111000000000000000000000011111110000000000111111111111110000000;
      map[64] = 160'b00000000001111111101111110000000111111101111111000000000000000000000000011111111000000000000000000000011111110000000001111111111111110000000;
      map[63] = 160'b00000000001111111001111110000000111111100111111000000000000000000000000011111111000000000000000000000011111110000000001111111011111110000000;
      map[62] = 160'b00000000001111111001111110000000111111100111111000000000000000000000000011111111000000000000000000000011111110000000011111110011111110000000;
      map[61] = 160'b00000000011111111001111110000001111111100111111100000000000000000000000011111111000000000000000000000011111110000000111111110011111110000000;
      map[60] = 160'b00000000011111111000111111000001111111000111111100000000000000000000000011111111000000000000000000000011111110000000111111100011111110000000;
      map[59] = 160'b00000000011111110000111111000001111111000011111100000000000000000000000011111111000000000000000000000011111110000001111111100011111110000000;
      map[58] = 160'b00000000011111110000111111000001111111000011111100000000000000000000000011111111000000000000000000000011111110000011111111000011111110000000;
      map[57] = 160'b00000000111111110000011111000011111111000011111110000000000000000000000011111111000000000000000000000011111110000011111110000011111110000000;
      map[56] = 160'b00000000111111110000011111100011111110000011111110000000000000000000000011111111000000000000000000000011111110000111111110000011111110000000;
      map[55] = 160'b00000000111111110000011111100011111110000011111110000000000000000000000011111111000000000000000000000011111110000111111100000011111110000000;
      map[54] = 160'b00000000111111100000011111100011111110000011111110000000000000000000000011111111000000000000000000000011111110001111111000000011111110000000;
      map[53] = 160'b00000001111111100000011111110111111110000011111110000000000000000000000011111111000000000000000000000011111110001111111000000011111110000000;
      map[52] = 160'b00000001111111100000011111110111111100000011111110000000000000000000000011111111000000000000000000000011111110001111111000000011111110000000;
      map[51] = 160'b00000001111111100000011111110111111100000011111110000000000000000000000011111111000000000000000000000011111110011111110000000011111110000000;
      map[50] = 160'b00000001111111000000001111110111111100000011111111000000000000000000000011111111000000000000000000000011111110111111110000000011111110000000;
      map[49] = 160'b00000001111111000000001111111111111100000001111111000000000000000000000011111111000000000000000000000011111110111111100000000011111110000000;
      map[48] = 160'b00000001111111000000001111111111111000000001111111000000000000000000000011111111000000000000000000000011111111111111000000000011111110000000;
      map[47] = 160'b00000001111111000000001111111111111000000001111111000000000000000000000011111111000000000000000000000011111111111111000000000011111110000000;
      map[46] = 160'b00000001111111000000000111111111111000000001111111100000000000000000000011111111000000000000000000000011111111111110000000000011111110000000;
      map[45] = 160'b00000011111111000000000111111111111000000001111111100000000000000000000011111111000000000000000000000011111111111110000000000011111110000000;
      map[44] = 160'b00000011111111000000000111111111111000000000111111100000000000000000000011111111000000000000000000000011111111111100000000000011111110000000;
      map[43] = 160'b00000011111111000000000111111111111000000000111111100000000000000000001111111111111000000000000000000011111111111000000000000011111110000000;
      map[42] = 160'b00000111111111000000000011111111111000000000111111110000000000000000001111111111111000000000000000000011111111111000000000000011111110000000;
      map[41] = 160'b00000111111110000000000011111111111000000000111111110000000000000000001111111111111000000000000000000011111111110000000000000011111110000000;
      map[40] = 160'b00000111111110000000000011111111110000000000011111110000000000000000001111111111111000000000000000000011111111110000000000000011111110000000;
      map[39] = 160'b00000111111110000000000001111111110000000000011111111000000000000000001111111111111000000000000000000011111111110000000000000011111110000000;
      map[38] = 160'b00001111111110000000000001111111110000000000011111111000000000000000001111111111111000000000000000000011111111100000000000000011111110000000;
      map[37] = 160'b00001111111110000000000001111111110000000000011111111000000000000000001111111111111000000000000000000011111111000000000000000011111110000000;
      map[36] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[35] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[34] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[33] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[32] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[31] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[30] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[29] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[28] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[27] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[26] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[25] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[24] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[23] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[22] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[21] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[20] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[19] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[18] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[17] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[16] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[15] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[14] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[13] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[12] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[11] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[10] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[9] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[8] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[7] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[6] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[5] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[4] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[3] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[2] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      map[1] = 160'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	end
//	clk1ms m4(clk, clk_1ms);
	always @(posedge clk) begin
		if (py>180 && py<=300 && px>240 && px<=400) out <= ((map[py-180] & (1<<(400-px)))>0) ? 1 : 0;
	end
	assign end_on = out;
endmodule
