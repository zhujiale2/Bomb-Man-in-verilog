`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:30:40 01/07/2014 
// Design Name: 
// Module Name:    bombmask 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bombmask(
	input wire clk,
	input wire [9:0] px, py,
	output wire [2:0] col
);
	reg [0:15] green [0:15];
	reg [0:15] blue [0:15];
	reg [0:15] red [0:15];
	initial begin
      green[15] = 16'b0000000000000000;
      green[14] = 16'b0000000000000000;
      green[13] = 16'b0000000000000000;
      green[12] = 16'b0000000000000000;
      green[11] = 16'b0000000000000000;
      green[10] = 16'b0000000000000000;
      green[9]  = 16'b0000000000000000;
      green[8]  = 16'b0000000000000000;
      green[7]  = 16'b0000100000000000;
      green[6]  = 16'b0000100000000000;
      green[5]  = 16'b0000011000000000;
      green[4]  = 16'b0000001100000000;
      green[3]  = 16'b0000000000000000;
      green[2]  = 16'b0000000000000000;
      green[1]  = 16'b0000000000000000;
      green[0]  = 16'b0000000000000000;
		
		
		
		blue[15] = 16'b0000000000000000;
      blue[14] = 16'b0000000000000000;
      blue[13] = 16'b0000000000000000;
      blue[12] = 16'b0000000000000000;
      blue[11] = 16'b0000000000000000;
      blue[10] = 16'b0000000000000000;
      blue[9]  = 16'b0000000000000000;
      blue[8]  = 16'b0000000000000000;
      blue[7]  = 16'b0000100000000000;
      blue[6]  = 16'b0000100000000000;
      blue[5]  = 16'b0000011000000000;
      blue[4]  = 16'b0000001100000000;
      blue[3]  = 16'b0000000000000000;
      blue[2]  = 16'b0000000000000000;
      blue[1]  = 16'b0000000000000000;
      blue[0]  = 16'b0000000000000000;
		
		red[15] = 16'b0000001111000000;
      red[14] = 16'b0000110000110000;
      red[13] = 16'b0011100000011100;
      red[12] = 16'b0010000000000100;
      red[11] = 16'b0110000000000110;
      red[10] = 16'b0100000000000010;
      red[9]  = 16'b1000000000000001;
      red[8]  = 16'b1000000000000001;
      red[7]  = 16'b1000100000000001;
      red[6]  = 16'b1000100000000001;
      red[5]  = 16'b0100011000000010;
      red[4]  = 16'b0110001100000110;
      red[3]  = 16'b0010000000000100;
      red[2]  = 16'b0011100000011100;
      red[1]  = 16'b0000110000110000;
      red[0]  = 16'b0000001111000000;
	end
	assign col[2] = (green[py%16] & (1<<(15-px%16)))>0 ? 1 : 0;
	assign col[1] = (blue[py%16] & (1<<(15-px%16)))>0 ? 1 : 0;
	assign col[0] = (red[py%16] & (1<<(15-px%16)))>0 ? 1 : 0;
endmodule
