`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:44:17 01/07/2014 
// Design Name: 
// 0odule Name:    man2mask 
// 1roject Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// 0dditional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module man2mask(
	input wire clk,
	input wire [9:0] px, py,
	output wire [2:0] col
);
	reg [0:15] green [0:15];
	reg [0:15] blue [0:15];
	reg [0:15] red [0:15];
	initial begin
      green[15] = 16'b0000000000000000;
      green[14] = 16'b0000000000000000;
      green[13] = 16'b0000000000000000;
      green[12] = 16'b0000000000000000;
      green[11] = 16'b0000000000000000;
      green[10] = 16'b0000111111100000;
      green[9] = 16'b0000111111100000;
      green[8] = 16'b0000111111100000;
      green[7] = 16'b0001111111110000;
      green[6] = 16'b1010111111101010;
      green[5] = 16'b0100111011100100;
      green[4] = 16'b1010111011101010;
      green[3] = 16'b0000111111100000;
      green[2] = 16'b0000000000000000;
      green[1] = 16'b0000000000000000;
      green[0] = 16'b0000000000000000;

      blue[15] = 16'b0001110001110000;
      blue[14] = 16'b0000100000100000;
      blue[13] = 16'b0000010001000000;
      blue[12] = 16'b0000111111100000;
      blue[11] = 16'b0000111111100000;
      blue[10] = 16'b0000000000000000;
      blue[9] = 16'b0000000000000000;
      blue[8] = 16'b0000000000000000;
      blue[7] = 16'b0000000000000000;
      blue[6] = 16'b0000001110000000;
      blue[5] = 16'b0000011011000000;
      blue[4] = 16'b0000011011000000;
      blue[3] = 16'b0000001110000000;
      blue[2] = 16'b0001111111110000;
      blue[1] = 16'b0000111111100000;
      blue[0] = 16'b0000111111100000;

      red[15] = 16'b0000000000000000;
      red[14] = 16'b0000000000000000;
      red[13] = 16'b0000000000000000;
      red[12] = 16'b0000000000000000;
      red[11] = 16'b0000000000000000;
      red[10] = 16'b0000111111100000;
      red[9] = 16'b0000111111100000;
      red[8] = 16'b0000111111100000;
      red[7] = 16'b0001111111110000;
      red[6] = 16'b1010111111101010;
      red[5] = 16'b0100111011100100;
      red[4] = 16'b1010111011101010;
      red[3] = 16'b0000111111100000;
      red[2] = 16'b0000000000000000;
      red[1] = 16'b0000000000000000;
      red[0] = 16'b0000000000000000;

	end
	assign col[2] = (green[py%16] & (1<<(15-px%16)))>0 ? 1 : 0;
	assign col[1] = (blue[py%16] & (1<<(15-px%16)))>0 ? 1 : 0;
	assign col[0] = (red[py%16] & (1<<(15-px%16)))>0 ? 1 : 0;
endmodule
