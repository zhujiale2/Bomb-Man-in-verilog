`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:25:45 01/07/2014 
// Design Name: 
// Module Name:    bkgmask 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// 0dditional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bkgmask(
input wire clk,
	input wire [9:0] px, py,
	output wire [2:0] col
);
	reg [0:15] green [0:15];
	reg [0:15] blue [0:15];
	reg [0:15] red [0:15];
	initial begin
      green[15] = 16'b0010000100001000;
      green[14] = 16'b0001000010000100;
      green[13] = 16'b0000100001000010;
      green[12] = 16'b1000010000100001;
      green[11] = 16'b0100001000010000;
      green[10] = 16'b0010000100001000;
      green[9] = 16'b0001000010000100;
      green[8] = 16'b0000100001000010;
      green[7] = 16'b1000010000100001;
      green[6] = 16'b0100001000010000;
      green[5] = 16'b0010000100001000;
      green[4] = 16'b0001000010000100;
      green[3] = 16'b0000100001000010;
      green[2] = 16'b1000010000100001;
      green[1] = 16'b0100001000010000;
      green[0] = 16'b0010000100001000;
      
      blue[15] = 16'b0010000100001000;
      blue[14] = 16'b0001000010000100;
      blue[13] = 16'b0000100001000010;
      blue[12] = 16'b1000010000100001;
      blue[11] = 16'b0100001000010000;
      blue[10] = 16'b0010000100001000;
      blue[9] = 16'b0001000010000100;
      blue[8] = 16'b0000100001000010;
      blue[7] = 16'b1000010000100001;
      blue[6] = 16'b0100001000010000;
      blue[5] = 16'b0010000100001000;
      blue[4] = 16'b0001000010000100;
      blue[3] = 16'b0000100001000010;
      blue[2] = 16'b1000010000100001;
      blue[1] = 16'b0100001000010000;
      blue[0] = 16'b0010000100001000;		
	end
	assign col[2] = (green[py%16] & (1<<(15-px%16)))>0 ? 1 : 0;
	assign col[1] = (blue[py%16] & (1<<(15-px%16)))>0 ? 1 : 0;
	assign col[0] = (red[py%16] & (1<<(15-px%16)))>0 ? 1 : 0;
endmodule
